module ControlUnit(input [5:0]opcode, output RegDst, output Branch, output MemRead, output MemtoReg, 
						output ALUOp, output MemWrite, output ALUSrc, output RegWrite);
//	
//	always @(opcode)
//		begin 
//		case(<opcode>)
//			if ()
//		end
endmodule