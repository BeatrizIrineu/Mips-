module ArithmeticLogicUnit(input [31:0]readData1, input [31:0]readData2, input ALUControl);


endmodule 