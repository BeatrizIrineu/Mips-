module signExtend #(parameter N=31)
						(input [15:0] case1, input [25:0] case2, input [31:0] case3, output [N:0] sign_extended);

//  assign extended_value = {{16{input_value[15]}}, input_value};

 endmodule
