module ArithmeticLogicUnit(input [0:31]readData1, input [0:31]readData2, input ALUControl);


endmodule 